module alu_tb;
    reg     [5:0]   A, B;	// 測試輸入操作數 A 和 B，6 位元
	reg		[3:0]	op;		// 測試輸入操作碼，4 位元
    wire    [5:0]   Y;		// 測試輸出結果，6 位元

    // 實例化 ALU 模組，名稱為 m0，連接測試輸入和輸出
	alu m0(A, B, op, Y);
	
    // 使用 $monitor 顯示模擬時間和變數值
	initial
		$monitor("Time: %3t ns, A = %6b, B = %6b, op = %4b, Y = %6b", 
		         $time, A, B, op, Y);

	initial begin
        // 第一組測試案例：A = 13, B = 7，測試所有運算操作碼
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h0; // 測試操作碼 0
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h1; // 測試操作碼 1
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h2; // 測試操作碼 2
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h3; // 測試操作碼 3
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h4; // 測試操作碼 4
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h5; // 測試操作碼 5
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h6; // 測試操作碼 6
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h7; // 測試操作碼 7
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h8; // 測試操作碼 8
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'h9; // 測試操作碼 9
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'hA; // 測試操作碼 A
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'hB; // 測試操作碼 B
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'hC; // 測試操作碼 C
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'hD; // 測試操作碼 D
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'hE; // 測試操作碼 E
        #10 A = 6'd13; 	B = 6'd7; 	op = 4'hF; // 測試操作碼 F
		
		// 第二組測試案例：A = 5, B = 12，測試所有運算操作碼
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h0; // 測試操作碼 0
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h1; // 測試操作碼 1
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h2; // 測試操作碼 2
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h3; // 測試操作碼 3
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h4; // 測試操作碼 4
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h5; // 測試操作碼 5
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h6; // 測試操作碼 6
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h7; // 測試操作碼 7
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h8; // 測試操作碼 8
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'h9; // 測試操作碼 9
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'hA; // 測試操作碼 A
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'hB; // 測試操作碼 B
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'hC; // 測試操作碼 C
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'hD; // 測試操作碼 D
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'hE; // 測試操作碼 E
        #10 A = 6'd5; 	B = 6'd12; 	op = 4'hF; // 測試操作碼 F
        
		// 模擬結束
		#20 $finish;
	end
endmodule